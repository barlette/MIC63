.SUBCKT PASS GND IN OUT VDD
MM0 VDD IN OUT VDD pmos_rvt w=81n l=20n nfin=3
MM1 VDD IN OUT VDD pmos_rvt w=81n l=20n nfin=3
MM2 OUT IN GND GND nmos_rvt w=81n l=20n nfin=3
MM3 OUT IN GND GND nmos_rvt w=81n l=20n nfin=3
.ENDS
